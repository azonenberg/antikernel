localparam TX_SYMBOL_N2			= 0;	//-2.5V
localparam TX_SYMBOL_N1			= 1;	//-1V
localparam TX_SYMBOL_0			= 2;	// 0V
localparam TX_SYMBOL_1			= 3;	//+1V
localparam TX_SYMBOL_2			= 4;	//+2.5V
